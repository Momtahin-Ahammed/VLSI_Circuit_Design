// DSCH 3.5
// 15-Mar-22 11:40:50 PM
// E:\SPRING 2022\VLSI\LAB\ALU_drawing.sch

module ALU_drawing( );
endmodule

// Simulation parameters in Verilog Format

// Simulation parameters
